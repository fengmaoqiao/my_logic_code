// *********************************************************************************
// Project Name :
// Author       : libing
// Email        : lb891004@163.com
// Creat Time   : 2014/2/18 17:11:55
// File Name    : uart_driver.v
// Module Name  : uart_driver
// Called By    : 
// Abstract     :
//
// CopyRight(c) 2014, Zhimingda digital equipment Co., Ltd.. 
// All Rights Reserved
//
// *********************************************************************************
// Modification History:
// 1. initial
// *********************************************************************************/
// *************************
// MODULE DEFINITION
//
// Hierarchy:
// uart_driver
//     |---> uart_send
//     |---> uart_receive
// *************************
`timescale 1 ns / 1 ps

module uart_debug_driver(
//-----------------------------------------------------------------------------------
//Global Sinals 
//-----------------------------------------------------------------------------------     
    input               rst_n                   ,   // Reset, Valid low  
    input               clk_uart                ,   // Uart Refence Clock  
    input               baud_en                 ,   // Baudrate Enable, Last 1 clock cycle  
//-----------------------------------------------------------------------------------
//Software Config Sinals 
//-----------------------------------------------------------------------------------  
    input               verify_en               ,   // Verify Enable, 1-Enable; 0-Disable
    input               verify_select           ,   // Verify Mode Select, 1-Odd; 0-Even
    input               stop_bit_sel            ,   // Stop Bit Width Select, 1-2 bit; 0-1 bit 
    input               verify_filter           ,   // Verify faild filter,  1-Enable; 0-Disable
    input [3:0]         data_width              ,   // Data Width, valid rang: 8~5
//-----------------------------------------------------------------------------------
//Tx Data Load Interface
//-----------------------------------------------------------------------------------                                                   
    input [7:0]         tx_data                 ,   // TX data
    input               tx_start                ,   // TX start signal, Valid high
//-----------------------------------------------------------------------------------
//Rx data Sinals 
//-----------------------------------------------------------------------------------    
    output [7:0]        rx_data                 ,   // Recieved Data  
    output              rx_data_vld             ,   // Recieved Data Strobe, Last 1 baudrate cycle    
//-----------------------------------------------------------------------------------
//Software Interface Sinals 
//-----------------------------------------------------------------------------------     
    output              tx_busy                 ,   // TX busy, 1-busy; 0-idle
//-----------------------------------------------------------------------------------
//TX-Line & RX-Line Sinals
//-----------------------------------------------------------------------------------     
    input               rx_in                   ,   // UART Recieve Line
    output              tx_out                      // UART Transmit Line  
);


uart_debug_receive u_uart_receive(
//-----------------------------------------------------------------------------------
//Global Sinals 
//-----------------------------------------------------------------------------------     
    .rst_n                      (rst_n                      ),
    .clk_uart                   (clk_uart                   ),
    .baud_en                    (baud_en                    ),
//-----------------------------------------------------------------------------------
//Software Interface Sinals 
//-----------------------------------------------------------------------------------   
    .verify_en                  (verify_en                  ),
    .verify_select              (verify_select              ),
    .verify_filter              (verify_filter              ),
    .data_width                 (data_width                 ),
//-----------------------------------------------------------------------------------
//RX-Line Sinals
//----------------------------------------------------------------------------------- 
    .rx_in                      (rx_in                      ),
//-----------------------------------------------------------------------------------
//Rx data Sinals 
//-----------------------------------------------------------------------------------    
    .rx_data                    (rx_data                    ),
    .rx_data_vld                (rx_data_vld                )
);


uart_debug_send u_uart_send(
//-----------------------------------------------------------------------------------
//Global Sinals 
//-----------------------------------------------------------------------------------     
    .rst_n                      (rst_n                      ),
    .clk_uart                   (clk_uart                   ),
    .baud_en                    (baud_en                    ),
//-----------------------------------------------------------------------------------
//Software Config Sinals 
//-----------------------------------------------------------------------------------  
    .verify_en                  (verify_en                  ),
    .verify_select              (verify_select              ),
    .stop_bit_sel               (stop_bit_sel               ),
    .data_width                 (data_width                 ),
//-----------------------------------------------------------------------------------
//Tx Data Load Interface
//-----------------------------------------------------------------------------------                                                   
    .tx_data                    (tx_data                    ),
    .tx_start                   (tx_start                   ),
//-----------------------------------------------------------------------------------
//Software Interface Sinals 
//-----------------------------------------------------------------------------------     
    .tx_busy                    (tx_busy                    ),
//-----------------------------------------------------------------------------------
//TX-Line Sinals
//-----------------------------------------------------------------------------------     
    .tx_out                     (tx_out                     )
);


endmodule





